Blue
0 0 0 0 0 h 1 B 9 B 
0 0 0 0 0 h 3 B 11 B 
0 0 0 0 0 h 5 B 19 B 
0 0 0 0 0 h 7 B 21 B 
0 11 2 8 4 3 0 10 3 9 2 6 1 5 1 3 3 8 2 12 0 11 3 5 1 4 0 4 1 6 4 10 4 2 5 7 2 9 
17
